circuito de controle de ganho - chave

*-----------------------------Cabecalho-----------------------------*
*Criador: Gustavo Pinheiro
*email: gustavo.pinheiro@ufabc.edu.br
*data: 11/2024
*objetivo: Verificar o funcionamento do circuito de controle de ganho com uso de chave digital.
* O sinal a ser amplificado eh conectado a um Amplificador não-inversor, com o resistor de
*feedback sendo "Rf". Ja o resistor Rs num conjunto de resistores em paralelo, para controlar o ganho da saida.
*-------------------------------------------------------------------------------*

*----------------------Descricao dos modelos utilizados-------------------------*
* Comando incluir o conteúdo do subcircuito do AD826A:
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
*.SUBCKT AD826A  2  1  99 50 46
.include ad826a.cir

*.model diode_model D
.include 1N4148.cir;           diodo de pequenos sinais
*-------------------------------------------------------------------------------*


*-----------------------------Descricao do circuito-----------------------------*
*.param A=0.3 f=250k T={1/f}

*vSinal  vin     GND     sin(0 A f)
vSinal  vin     GND     AC 0.5V
VCC     vcc     GND     9V
VEE     vee     GND     -9V
*Cx      no2     no1      100n
*Rx      no2     GND     510
X_U1    vin     no1     vcc     vee     no1     AD826A
X_U2    GND     vrh     vcc     vee     out     AD826A
Rin     vrh     no1     1k


R0      tmp1    vrh      300
*R1      tmp2    tmp1     620
*R2      tmp3    tmp2     1.3k
R3      tmp4    tmp3     5.1k
*R4      out     tmp4     10k

C1      tmp1    GND    5p
C2      tmp2    GND    5p
C3      tmp3    GND    5p
C4      tmp4    GND    5p

*Raux1   tmp2    tmp1    180 ; resistores auxiliares Raux, para corrigir o erro "Singular matrix warning", gerado por
*Raux2   tmp3    tmp2    180   ; um nó de impedância infinita (por exemplo, uma conexão em série de dois capacitores)
Raux3   tmp4    tmp3    180      ;https://electronics.stackexchange.com/questions/361906/singular-matrix-warning
*Raux4   out     tmp4    180



Rcarga  out     GND     1k


*-------------------------------------------------------------------------------*


*-----------------------------Parametros de simulacao----------------------------*
.ac     dec     100     100     10Mega
*-------------------------------------------------------------------------------*

*-----------------------------Parametros de output----------------------------*
.control
    destroy all
    run
    plot vin out
    plot vin db(out-vin)
.endc

*-------------------------------------------------------------------------------*

.end
