Fonte de corrente com controle automatico de ganho

*-----------------------------Cabecalho-----------------------------*
*Criador: Gustavo Pinheiro
*email: gustavo.pinheiro@ufabc.edu.br
*data: 03/2024
*objetivo: Realizar o controle do ganho de uma fonte de corrente howland aperfeicoada por meio do 
*potenciometro digital. 
*A saida da fonte de corrente eh conectada a um Amplificador não-inversor, com o resistor de 
*feedback sendo "R2". Ja o resistor Rs varia entre 1k e 100k ohms, para controlar o ganho a saida vout
*-------------------------------------------------------------------------------*


*----------------------Descricao dos modelos utilizados-------------------------*
* Comando incluir o conteúdo do subcircuito do AD826A:
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
*.SUBCKT AD826A  2  1  99 50 46
.include ad826a.cir

*.model diode_model D
.include 1N4148.cir;           diodo de pequenos sinais
*-------------------------------------------------------------------------------*


*-----------------------------Descricao do circuito-----------------------------*
.param A=1 f=250k T={1/f}

vSinal	vin	GND	sin(0 A f)
VCC     vcc     GND     9V
VEE     vee     GND     -9V
C1	vin	v1	1.6u
R1	v1	GND	10k
X_U1	v1	v2	vcc	vee	v2	AD826A
X_U2	v2	vrh	vcc	vee	vout	AD826A
R2	vout	vrh	100k
Rs	vrh	GND	1k

C1b	vout	vout2	1.6u
R1b	vout2	GND	10k
*-------------------------------------------------------------------------------*



*-----------------------------Parametros de simulacao----------------------------*
*.ac	dec	100	100	10Mega
.tran {T/10000} {5*T}; simulacao transiente, 10000 passos por periodo, por 1,1 periodo
*-------------------------------------------------------------------------------*



*-----------------------------Parametros de output----------------------------*
.control
	let start_r = 10k
	let stop_r  = 100k
	let delta_r = {stop_r/10} ;{stop_r/num de simulacoes}

 	 let r_act = start_r
	 while r_act le stop_r ;realiza uma simulacao transciente (.tran) para cada passo de Rs
    		alter Rs r_act
    		run
    		let r_act = r_act + delta_r
  	end

set plotstyle=linplot;                  Retorna ao estilo default de plotagem
set color0=white;                       Muda a cor do background
set color1=black;                        Muda a cor da borda e do grid
set xbrushwidth=1; ; espessura das linhas
set hcopypscolor=1 ; para deixar arquivo .ps colorido

foreach iter 1 2 3 4 5 6 7 8 9 10 			; 10 simulacoes realizadas
*foreach iter 6 7 8 9 10				; ou escolher x (nesse exemplo sao 5) simulacoes entre as 10 realizadas
	let sim_{$iter} = tran{$iter}.v(vout)		; salva o sinal de saída para cada simulacao .tran
		meas tran atraso{$iter}		; calcula o atraso entre cada saida e a entrada
		+ TRIG v(vin)	VAL=0	FALL=1 TARG V(sim_{$iter}) VAL=0	FALL=1
end

plot vin sim_1 sim_2 sim_3 Sim_4 sim_5 	; plota as 5 primeiras simulacoes 
    hardcopy fonte_1.ps  vin sim_1 sim_2 sim_3 Sim_4 sim_5  
plot vin sim_6 sim_7 sim_8 Sim_9 sim_10 	; plota as 5 ultimas simulacoes
    hardcopy fonte_corrente_2.ps  vin sim_6 sim_7 sim_8 Sim_9 sim_10   

*----atraso do sinal
foreach iter 1 2 3 4 5 6 7 8 9 10 
	print  atraso{$iter}*180*2*250k 	;atraso do sinal para cada simulacao, em graus
end

let grau = 180*2*250k
plot atraso1*grau atraso2*grau atraso3*grau atraso4*grau atraso5*grau
+ atraso6*grau atraso7*grau atraso8*grau atraso9*grau atraso10*grau		;imprime os atrasos
    hardcopy fonte_corrente_atraso.ps  atraso1*grau atraso2*grau atraso3*grau atraso4*grau atraso5*grau   
    +atraso6*grau atraso7*grau atraso8*grau atraso9*grau atraso10*grau	
    
.endc
*-------------------------------------------------------------------------------*
.end
